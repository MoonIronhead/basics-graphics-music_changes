// Board configuration: tang_nano_9k_lcd_480_272_tm1638_hackathon
// This module uses few parameterization and relaxed typing rules

module hackathon_top
(
    input  logic       clock,
    input  logic       slow_clock,
    input  logic       reset,

    input  logic [7:0] key,
    output logic [7:0] led,

    // A dynamic seven-segment display

    output logic [7:0] abcdefgh,
    output logic [7:0] digit,

    // LCD screen interface

    input  logic [8:0] x,
    input  logic [8:0] y,

    output logic [4:0] red,
    output logic [5:0] green,
    output logic [4:0] blue
);

    always_comb
    begin
        red   = 0;
        green = 0;
        blue  = 0;

        if (x > 100 & x < 300 & y > 50 & y < 100)
            red = 31;

        // 31 is the maximum 5-bit number, 5'b11111

        // Exercise 1: Uncomment the code for a green rectangle
        // that overlaps red rectangle

        if (key[0])
        begin
            if (x > 200 & x < 400 & y > 150 & y < 200)
            green = 63;
        end
        else
        begin
            if (x > 120 & x < 320 & y > 70 & y < 120)
            blue = 63;
        end

        // 63 is the maximum 6-bit number, 6'b111111

        // Excersice 2: Make a circle

        begin
            int radius = 50;
            int center_x = 240;
            int center_y = 136;

            if ((x - center_x) * (x - center_x) + (y - center_y) * (y - center_y) <= radius*radius)
                blue = 63;
        end

        // Exercise 2: Add a blue rectangle
        // that overlaps both rectangles

        if (x > 150 & x < 250 & y > 100 & y < 150)
            blue = 31;

    end
endmodule
